** sch_path: /home/ttuser/tt06-OTA-Simmettrico/xschem/Polarizzazione0.sch
**.subckt Polarizzazione0
Vgs net1 GND 0
Vds net2 GND 1.8
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice




 this option enables mos model bin
* selection based on W/NF instead of W
.opton wnflag=1
.option savecurrents


dc Vgs 0 1.8 0.2


set appendwrite
op

.end




**** end user architecture code
**.ends
.GLOBAL GND
.end
