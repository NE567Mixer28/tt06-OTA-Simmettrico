** sch_path: /home/ttuser/tt06-OTA-Simmettrico/xschem/Polarizzazione0.sch
**.subckt Polarizzazione0
Vgs GND net1 1
Vds GND net2 1.8
XM1 net3 net1 GND GND sky130_fd_pr__pfet_01v8_hvt L=1 W=Wp nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas net3 net2 0
.save i(vmeas)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice




.control
.param Wp =6
dc Vds 0 1.8 0.02 Vgs 0 1.4 0.2
 *let start_w = 1
  *let stop_w = 90
  *let delta_w = 5
  *let w_act = start_w
  *while w_act le stop_w
   * alterparam Wp = $&w_act
    *reset
   * save all
    *run
    *remzerovec
    *let w_act = w_act + delta_w
    plot i(Vds)
plot i(Vmeas)
write Polarizzazione0.raw


.endc
.save all




**** end user architecture code
**.ends
.GLOBAL GND
.end
