** sch_path: /home/ttuser/tt06-OTA-Simmettrico/xschem/Polarizzazione.sch
**.subckt Polarizzazione
XM2 vds vgs GND GND sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vgs GND vgs 0
vds GND vds 0
**** begin user architecture code


.dc vgs 0 1.8 1m vds 0 1.8  1m
.save all
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
