** sch_path: /home/ttuser/tt06-OTA-Simmettrico/xschem/Polarizzazione.sch
**.subckt Polarizzazione
XM2 net1 Vbias GND VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 GND Vbias 1
V2 GND net1 1.8
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.op



**** end user architecture code
**.ends
.GLOBAL GND
.end
